magic
tech sky130A
magscale 1 2
timestamp 1745678094
<< checkpaint >>
rect -3932 -3108 10832 14396
<< viali >>
rect 4997 9129 5031 9163
rect 5365 9061 5399 9095
rect 1409 8993 1443 9027
rect 1685 8925 1719 8959
rect 2329 8925 2363 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 2513 8789 2547 8823
rect 1777 8449 1811 8483
rect 4905 8449 4939 8483
rect 5181 8449 5215 8483
rect 1869 8381 1903 8415
rect 2145 8381 2179 8415
rect 4997 8381 5031 8415
rect 4905 8245 4939 8279
rect 5365 8245 5399 8279
rect 1593 8041 1627 8075
rect 2513 8041 2547 8075
rect 1409 7837 1443 7871
rect 2329 7837 2363 7871
rect 5181 7837 5215 7871
rect 5365 7701 5399 7735
rect 1409 7361 1443 7395
rect 1501 7361 1535 7395
rect 3893 7361 3927 7395
rect 4169 7361 4203 7395
rect 1685 7293 1719 7327
rect 3985 7293 4019 7327
rect 4077 7225 4111 7259
rect 1593 7157 1627 7191
rect 4353 7157 4387 7191
rect 1409 6749 1443 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 5181 6749 5215 6783
rect 4077 6681 4111 6715
rect 1593 6613 1627 6647
rect 4629 6613 4663 6647
rect 5365 6613 5399 6647
rect 3433 5321 3467 5355
rect 4905 5321 4939 5355
rect 4813 5253 4847 5287
rect 1409 5185 1443 5219
rect 3249 5185 3283 5219
rect 4721 5185 4755 5219
rect 5181 5117 5215 5151
rect 1593 4981 1627 5015
rect 4077 4777 4111 4811
rect 5365 4777 5399 4811
rect 4261 4709 4295 4743
rect 3893 4641 3927 4675
rect 4629 4641 4663 4675
rect 5089 4641 5123 4675
rect 4077 4573 4111 4607
rect 4721 4573 4755 4607
rect 5181 4573 5215 4607
rect 3801 4505 3835 4539
rect 1869 4233 1903 4267
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 2605 4097 2639 4131
rect 4629 4097 4663 4131
rect 4905 4097 4939 4131
rect 4997 4097 5031 4131
rect 5181 4097 5215 4131
rect 2697 4029 2731 4063
rect 4721 4029 4755 4063
rect 4169 3961 4203 3995
rect 4353 3961 4387 3995
rect 1593 3893 1627 3927
rect 2605 3893 2639 3927
rect 2973 3893 3007 3927
rect 5365 3893 5399 3927
rect 3801 3689 3835 3723
rect 4169 3553 4203 3587
rect 3985 3485 4019 3519
rect 2053 3145 2087 3179
rect 1685 3009 1719 3043
rect 1777 2941 1811 2975
rect 1869 2601 1903 2635
rect 1593 2533 1627 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 1394 8984 1400 9036
rect 1452 8984 1458 9036
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 2332 8888 2360 8919
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 1268 8860 2360 8888
rect 1268 8848 1274 8860
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 5184 8888 5212 8919
rect 2464 8860 5212 8888
rect 2464 8848 2470 8860
rect 2498 8780 2504 8832
rect 2556 8780 2562 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 2498 8548 2504 8560
rect 1780 8520 2504 8548
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1780 8489 1808 8520
rect 2498 8508 2504 8520
rect 2556 8508 2562 8560
rect 1765 8483 1823 8489
rect 1765 8480 1777 8483
rect 1452 8452 1777 8480
rect 1452 8440 1458 8452
rect 1765 8449 1777 8452
rect 1811 8449 1823 8483
rect 2314 8480 2320 8492
rect 1765 8443 1823 8449
rect 2056 8452 2320 8480
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1728 8384 1869 8412
rect 1728 8372 1734 8384
rect 1857 8381 1869 8384
rect 1903 8412 1915 8415
rect 2056 8412 2084 8452
rect 2314 8440 2320 8452
rect 2372 8480 2378 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 2372 8452 4905 8480
rect 2372 8440 2378 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 5132 8452 5181 8480
rect 5132 8440 5138 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 1903 8384 2084 8412
rect 2133 8415 2191 8421
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2133 8381 2145 8415
rect 2179 8412 2191 8415
rect 2406 8412 2412 8424
rect 2179 8384 2412 8412
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 2498 8372 2504 8424
rect 2556 8412 2562 8424
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 2556 8384 4997 8412
rect 2556 8372 2562 8384
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 4893 8279 4951 8285
rect 4893 8276 4905 8279
rect 1636 8248 4905 8276
rect 1636 8236 1642 8248
rect 4893 8245 4905 8248
rect 4939 8245 4951 8279
rect 4893 8239 4951 8245
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5353 8279 5411 8285
rect 5353 8276 5365 8279
rect 5040 8248 5365 8276
rect 5040 8236 5046 8248
rect 5353 8245 5365 8248
rect 5399 8245 5411 8279
rect 5353 8239 5411 8245
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 1578 8032 1584 8084
rect 1636 8032 1642 8084
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 4798 8072 4804 8084
rect 2547 8044 4804 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4212 7840 5181 7868
rect 4212 7828 4218 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 2314 7392 2320 7404
rect 1535 7364 2320 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3844 7364 3893 7392
rect 3844 7352 3850 7364
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 4706 7392 4712 7404
rect 4203 7364 4712 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1636 7296 1685 7324
rect 1636 7284 1642 7296
rect 1673 7293 1685 7296
rect 1719 7324 1731 7327
rect 2498 7324 2504 7336
rect 1719 7296 2504 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4522 7324 4528 7336
rect 4019 7296 4528 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4522 7284 4528 7296
rect 4580 7324 4586 7336
rect 4982 7324 4988 7336
rect 4580 7296 4988 7324
rect 4580 7284 4586 7296
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 4062 7216 4068 7268
rect 4120 7216 4126 7268
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 3878 7188 3884 7200
rect 1627 7160 3884 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4614 7188 4620 7200
rect 4387 7160 4620 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 5074 6848 5080 6860
rect 1596 6820 5080 6848
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1596 6653 1624 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4430 6780 4436 6792
rect 4203 6752 4436 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 5166 6740 5172 6792
rect 5224 6740 5230 6792
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6712 4123 6715
rect 4982 6712 4988 6724
rect 4111 6684 4988 6712
rect 4111 6681 4123 6684
rect 4065 6675 4123 6681
rect 4982 6672 4988 6684
rect 5040 6672 5046 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4028 6616 4629 6644
rect 4028 6604 4034 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5352 3479 5355
rect 4154 5352 4160 5364
rect 3467 5324 4160 5352
rect 3467 5321 3479 5324
rect 3421 5315 3479 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5352 4951 5355
rect 5166 5352 5172 5364
rect 4939 5324 5172 5352
rect 4939 5321 4951 5324
rect 4893 5315 4951 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 4801 5287 4859 5293
rect 4801 5253 4813 5287
rect 4847 5284 4859 5287
rect 5074 5284 5080 5296
rect 4847 5256 5080 5284
rect 4847 5253 4859 5256
rect 4801 5247 4859 5253
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 3234 5176 3240 5228
rect 3292 5176 3298 5228
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4212 5188 4721 5216
rect 4212 5176 4218 5188
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 4890 5148 4896 5160
rect 4580 5120 4896 5148
rect 4580 5108 4586 5120
rect 4890 5108 4896 5120
rect 4948 5148 4954 5160
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4948 5120 5181 5148
rect 4948 5108 4954 5120
rect 5169 5117 5181 5120
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 4246 5012 4252 5024
rect 1627 4984 4252 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 4246 4972 4252 4984
rect 4304 5012 4310 5024
rect 4706 5012 4712 5024
rect 4304 4984 4712 5012
rect 4304 4972 4310 4984
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 4062 4768 4068 4820
rect 4120 4768 4126 4820
rect 5350 4768 5356 4820
rect 5408 4768 5414 4820
rect 4249 4743 4307 4749
rect 4249 4709 4261 4743
rect 4295 4709 4307 4743
rect 4249 4703 4307 4709
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 3844 4644 3893 4672
rect 3844 4632 3850 4644
rect 3881 4641 3893 4644
rect 3927 4641 3939 4675
rect 4264 4672 4292 4703
rect 4338 4672 4344 4684
rect 4264 4644 4344 4672
rect 3881 4635 3939 4641
rect 4338 4632 4344 4644
rect 4396 4672 4402 4684
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 4396 4644 4629 4672
rect 4396 4632 4402 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 5074 4632 5080 4684
rect 5132 4632 5138 4684
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4604 4123 4607
rect 4246 4604 4252 4616
rect 4111 4576 4252 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 5040 4576 5181 4604
rect 5040 4564 5046 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 3789 4539 3847 4545
rect 3789 4505 3801 4539
rect 3835 4536 3847 4539
rect 4890 4536 4896 4548
rect 3835 4508 4896 4536
rect 3835 4505 3847 4508
rect 3789 4499 3847 4505
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 1857 4267 1915 4273
rect 1857 4233 1869 4267
rect 1903 4264 1915 4267
rect 2958 4264 2964 4276
rect 1903 4236 2964 4264
rect 1903 4233 1915 4236
rect 1857 4227 1915 4233
rect 2958 4224 2964 4236
rect 3016 4264 3022 4276
rect 4062 4264 4068 4276
rect 3016 4236 4068 4264
rect 3016 4224 3022 4236
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 1596 4168 1808 4196
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1596 4128 1624 4168
rect 1443 4100 1624 4128
rect 1673 4131 1731 4137
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 842 4020 848 4072
rect 900 4060 906 4072
rect 1688 4060 1716 4091
rect 900 4032 1716 4060
rect 900 4020 906 4032
rect 1394 3952 1400 4004
rect 1452 3992 1458 4004
rect 1780 3992 1808 4168
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 4304 4168 5028 4196
rect 4304 4156 4310 4168
rect 2406 4088 2412 4140
rect 2464 4128 2470 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2464 4100 2605 4128
rect 2464 4088 2470 4100
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 4614 4088 4620 4140
rect 4672 4088 4678 4140
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 5000 4137 5028 4168
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 2685 4063 2743 4069
rect 2685 4060 2697 4063
rect 2556 4032 2697 4060
rect 2556 4020 2562 4032
rect 2685 4029 2697 4032
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 4430 4020 4436 4072
rect 4488 4060 4494 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4488 4032 4721 4060
rect 4488 4020 4494 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 1452 3964 1716 3992
rect 1780 3964 4169 3992
rect 1452 3952 1458 3964
rect 1578 3884 1584 3936
rect 1636 3884 1642 3936
rect 1688 3924 1716 3964
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 4338 3952 4344 4004
rect 4396 3952 4402 4004
rect 2593 3927 2651 3933
rect 2593 3924 2605 3927
rect 1688 3896 2605 3924
rect 2593 3893 2605 3896
rect 2639 3893 2651 3927
rect 2593 3887 2651 3893
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 4062 3924 4068 3936
rect 3007 3896 4068 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3292 3692 3801 3720
rect 3292 3680 3298 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 3789 3683 3847 3689
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 4614 3652 4620 3664
rect 1636 3624 4620 3652
rect 1636 3612 1642 3624
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 4154 3544 4160 3596
rect 4212 3544 4218 3596
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3936 3488 3985 3516
rect 3936 3476 3942 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 2041 3179 2099 3185
rect 2041 3145 2053 3179
rect 2087 3176 2099 3179
rect 5166 3176 5172 3188
rect 2087 3148 5172 3176
rect 2087 3145 2099 3148
rect 2041 3139 2099 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2958 3040 2964 3052
rect 1719 3012 2964 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 3970 2972 3976 2984
rect 1811 2944 3976 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 4706 2632 4712 2644
rect 1903 2604 4712 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 3786 2564 3792 2576
rect 1627 2536 3792 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 3786 2524 3792 2536
rect 3844 2524 3850 2576
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 1216 8848 1268 8900
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 2412 8848 2464 8900
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1400 8440 1452 8492
rect 2504 8508 2556 8560
rect 1676 8372 1728 8424
rect 2320 8440 2372 8492
rect 5080 8440 5132 8492
rect 2412 8372 2464 8424
rect 2504 8372 2556 8424
rect 1584 8236 1636 8288
rect 4988 8236 5040 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 4804 8032 4856 8084
rect 848 7828 900 7880
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 4160 7828 4212 7880
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2320 7352 2372 7404
rect 3792 7352 3844 7404
rect 4712 7352 4764 7404
rect 1584 7284 1636 7336
rect 2504 7284 2556 7336
rect 4528 7284 4580 7336
rect 4988 7284 5040 7336
rect 4068 7259 4120 7268
rect 4068 7225 4077 7259
rect 4077 7225 4111 7259
rect 4111 7225 4120 7259
rect 4068 7216 4120 7225
rect 3884 7148 3936 7200
rect 4620 7148 4672 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 848 6740 900 6792
rect 5080 6808 5132 6860
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4436 6740 4488 6792
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 4988 6672 5040 6724
rect 3976 6604 4028 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 4160 5312 4212 5364
rect 5172 5312 5224 5364
rect 5080 5244 5132 5296
rect 848 5176 900 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 4160 5176 4212 5228
rect 4528 5108 4580 5160
rect 4896 5108 4948 5160
rect 4252 4972 4304 5024
rect 4712 4972 4764 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 4068 4811 4120 4820
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 3792 4632 3844 4684
rect 4344 4632 4396 4684
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 4252 4564 4304 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 4988 4564 5040 4616
rect 4896 4496 4948 4548
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 2964 4224 3016 4276
rect 4068 4224 4120 4276
rect 848 4020 900 4072
rect 1400 3952 1452 4004
rect 4252 4156 4304 4208
rect 2412 4088 2464 4140
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 2504 4020 2556 4072
rect 4436 4020 4488 4072
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 4344 3995 4396 4004
rect 4344 3961 4353 3995
rect 4353 3961 4387 3995
rect 4387 3961 4396 3995
rect 4344 3952 4396 3961
rect 4068 3884 4120 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 3240 3680 3292 3732
rect 1584 3612 1636 3664
rect 4620 3612 4672 3664
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 3884 3476 3936 3528
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 5172 3136 5224 3188
rect 2964 3000 3016 3052
rect 3976 2932 4028 2984
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 4712 2592 4764 2644
rect 3792 2524 3844 2576
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 1214 9072 1270 9081
rect 1412 9042 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 1214 9007 1270 9016
rect 1400 9036 1452 9042
rect 1228 8906 1256 9007
rect 5354 9007 5410 9016
rect 1400 8978 1452 8984
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 1216 8900 1268 8906
rect 1216 8842 1268 8848
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 848 7880 900 7886
rect 846 7848 848 7857
rect 900 7848 902 7857
rect 846 7783 902 7792
rect 1412 7410 1440 8434
rect 1688 8430 1716 8910
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1596 8090 1624 8230
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 846 5128 902 5137
rect 846 5063 902 5072
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 860 3777 888 4014
rect 1412 4010 1440 7346
rect 1596 7342 1624 8026
rect 2332 7886 2360 8434
rect 2424 8430 2452 8842
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 8566 2544 8774
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2516 8430 2544 8502
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 4816 8090 4844 8910
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 2332 7410 2360 7822
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2332 6914 2360 7346
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2332 6886 2452 6914
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2424 4146 2452 6886
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2516 4078 2544 7278
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 1400 4004 1452 4010
rect 1400 3946 1452 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 846 3768 902 3777
rect 846 3703 902 3712
rect 1596 3670 1624 3878
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2976 3058 3004 4218
rect 3252 3738 3280 5170
rect 3804 4690 3832 7346
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3804 2582 3832 4626
rect 3896 3534 3924 7142
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 6662 4016 6734
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3988 2990 4016 6598
rect 4080 4826 4108 7210
rect 4172 5370 4200 7822
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4540 6798 4568 7278
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 4282 4108 4762
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4068 3936 4120 3942
rect 4172 3890 4200 5170
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 4622 4292 4966
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4214 4292 4558
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4356 4010 4384 4626
rect 4448 4078 4476 6734
rect 4540 5166 4568 6734
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4632 4146 4660 7142
rect 4724 6798 4752 7346
rect 5000 7342 5028 8230
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5092 6866 5120 8434
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4724 5030 4752 6734
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4120 3884 4200 3890
rect 4068 3878 4200 3884
rect 4080 3862 4200 3878
rect 4172 3602 4200 3862
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3792 2576 3844 2582
rect 3792 2518 3844 2524
rect 4632 2446 4660 3606
rect 4724 2650 4752 4558
rect 4908 4554 4936 5102
rect 5000 4622 5028 6666
rect 5092 5302 5120 6802
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 5370 5212 6734
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6361 5396 6598
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5368 4826 5396 4927
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4908 4146 4936 4490
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5092 2446 5120 4626
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5184 3194 5212 4082
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 1214 9016 1270 9072
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 846 7828 848 7848
rect 848 7828 900 7848
rect 900 7828 902 7848
rect 846 7792 902 7828
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 846 6432 902 6488
rect 846 5072 902 5128
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 846 3712 902 3768
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4936 5410 4992
rect 5354 3576 5410 3632
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 1209 9074 1275 9077
rect 0 9072 1275 9074
rect 0 9016 1214 9072
rect 1270 9016 1275 9072
rect 0 9014 1275 9016
rect 0 8984 800 9014
rect 1209 9011 1275 9014
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7850 907 7853
rect 798 7848 907 7850
rect 798 7792 846 7848
rect 902 7792 907 7848
rect 798 7787 907 7792
rect 798 7744 858 7787
rect 0 7654 858 7744
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 0 7624 800 7654
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__or4_2  _09_
timestamp 0
transform 1 0 4876 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_
timestamp 0
transform -1 0 5152 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_
timestamp 0
transform -1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _13_
timestamp 0
transform 1 0 1472 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _14_
timestamp 0
transform -1 0 4416 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _15_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _16_
timestamp 0
transform -1 0 4692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 0
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _18_
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp 0
transform 1 0 1564 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _20_
timestamp 0
transform 1 0 2576 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _21_
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform -1 0 4232 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform -1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _24_
timestamp 0
transform -1 0 5244 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 0
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_11
timestamp 0
transform 1 0 2116 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_23
timestamp 0
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_35
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_47
timestamp 0
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_34
timestamp 0
transform 1 0 4232 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_46
timestamp 0
transform 1 0 5336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_9
timestamp 0
transform 1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_21
timestamp 0
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_35
timestamp 0
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_18
timestamp 0
transform 1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_22
timestamp 0
transform 1 0 3128 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_26
timestamp 0
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_38
timestamp 0
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_45
timestamp 0
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 0
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 0
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 0
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_34
timestamp 0
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_40
timestamp 0
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_7
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_19
timestamp 0
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_36
timestamp 0
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_12
timestamp 0
transform 1 0 2208 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_16
timestamp 0
transform 1 0 2576 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_12
timestamp 0
transform 1 0 2208 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_24
timestamp 0
transform 1 0 3312 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_36
timestamp 0
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_40
timestamp 0
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_16
timestamp 0
transform 1 0 2576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal1 s 4876 5134 4876 5134 4 _00_
rlabel metal2 s 4002 4862 4002 4862 4 _01_
rlabel metal1 s 4600 4046 4600 4046 4 _02_
rlabel metal1 s 4508 7174 4508 7174 4 _03_
rlabel metal1 s 4278 4692 4278 4692 4 _04_
rlabel metal1 s 1518 4114 1518 4114 4 _05_
rlabel metal2 s 4186 4386 4186 4386 4 _06_
rlabel metal1 s 3956 3502 3956 3502 4 _07_
rlabel metal1 s 3542 3706 3542 3706 4 _08_
rlabel metal3 s 1050 10404 1050 10404 4 in[0]
rlabel metal3 s 958 9044 958 9044 4 in[1]
rlabel metal3 s 0 7624 800 7744 4 in[2]
port 5 nsew
rlabel metal3 s 0 6264 800 6384 4 in[3]
port 6 nsew
rlabel metal3 s 0 4904 800 5024 4 in[4]
port 7 nsew
rlabel metal3 s 0 3544 800 3664 4 in[5]
port 8 nsew
rlabel metal3 s 0 2184 800 2304 4 in[6]
port 9 nsew
rlabel metal3 s 1188 884 1188 884 4 in[7]
rlabel metal1 s 2530 4114 2530 4114 4 net1
rlabel metal1 s 2300 8398 2300 8398 4 net10
rlabel metal1 s 3818 5338 3818 5338 4 net11
rlabel metal1 s 5060 5338 5060 5338 4 net12
rlabel metal1 s 5106 4590 5106 4590 4 net13
rlabel metal1 s 3634 3162 3634 3162 4 net14
rlabel metal2 s 4646 3026 4646 3026 4 net15
rlabel metal2 s 5106 3536 5106 3536 4 net16
rlabel metal1 s 1564 3978 1564 3978 4 net2
rlabel metal1 s 2622 4046 2622 4046 4 net3
rlabel metal1 s 3358 6834 3358 6834 4 net4
rlabel metal1 s 4186 4590 4186 4590 4 net5
rlabel metal2 s 2990 4250 2990 4250 4 net6
rlabel metal1 s 3864 4658 3864 4658 4 net7
rlabel metal1 s 3312 2618 3312 2618 4 net8
rlabel metal1 s 3680 8058 3680 8058 4 net9
rlabel metal2 s 5014 9775 5014 9775 4 out[0]
rlabel metal3 s 5382 9061 5382 9061 4 out[1]
rlabel metal3 s 5382 7701 5382 7701 4 out[2]
rlabel metal2 s 5382 6477 5382 6477 4 out[3]
rlabel metal2 s 5382 4879 5382 4879 4 out[4]
rlabel metal2 s 5382 3757 5382 3757 4 out[5]
rlabel metal3 s 4830 2261 4830 2261 4 out[6]
rlabel metal2 s 5474 1615 5474 1615 4 out[7]
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 10344 800 10464 0 FreeSans 600 0 0 0 in[0]
port 3 nsew
flabel metal3 s 0 8984 800 9104 0 FreeSans 600 0 0 0 in[1]
port 4 nsew
flabel metal3 s 400 7684 400 7684 0 FreeSans 600 0 0 0 in[2]
flabel metal3 s 400 6324 400 6324 0 FreeSans 600 0 0 0 in[3]
flabel metal3 s 400 4964 400 4964 0 FreeSans 600 0 0 0 in[4]
flabel metal3 s 400 3604 400 3604 0 FreeSans 600 0 0 0 in[5]
flabel metal3 s 400 2244 400 2244 0 FreeSans 600 0 0 0 in[6]
flabel metal3 s 0 824 800 944 0 FreeSans 600 0 0 0 in[7]
port 10 nsew
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 600 0 0 0 out[0]
port 11 nsew
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 600 0 0 0 out[2]
port 13 nsew
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 600 0 0 0 out[3]
port 14 nsew
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 600 0 0 0 out[4]
port 15 nsew
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 600 0 0 0 out[5]
port 16 nsew
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 6100 824 6900 944 0 FreeSans 600 0 0 0 out[7]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
