magic
tech sky130A
magscale 1 2
timestamp 1745676085
<< viali >>
rect 4997 9129 5031 9163
rect 5365 9061 5399 9095
rect 1409 8993 1443 9027
rect 1685 8925 1719 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 1409 8449 1443 8483
rect 3157 8449 3191 8483
rect 3341 8449 3375 8483
rect 1593 8313 1627 8347
rect 3341 8313 3375 8347
rect 1409 7837 1443 7871
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 5181 7837 5215 7871
rect 1593 7701 1627 7735
rect 2697 7701 2731 7735
rect 5365 7701 5399 7735
rect 3065 7361 3099 7395
rect 4077 7361 4111 7395
rect 3157 7293 3191 7327
rect 3985 7293 4019 7327
rect 3433 7225 3467 7259
rect 4445 7157 4479 7191
rect 1409 6749 1443 6783
rect 4813 6749 4847 6783
rect 5273 6749 5307 6783
rect 5181 6681 5215 6715
rect 1593 6613 1627 6647
rect 5089 6613 5123 6647
rect 2973 6409 3007 6443
rect 5365 6409 5399 6443
rect 3249 6273 3283 6307
rect 5181 6273 5215 6307
rect 2973 6205 3007 6239
rect 3157 6069 3191 6103
rect 3525 5321 3559 5355
rect 4537 5321 4571 5355
rect 1685 5253 1719 5287
rect 1409 5185 1443 5219
rect 1961 5185 1995 5219
rect 2421 5185 2455 5219
rect 2697 5185 2731 5219
rect 3157 5185 3191 5219
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 1777 5117 1811 5151
rect 2513 5117 2547 5151
rect 3065 5117 3099 5151
rect 4077 5117 4111 5151
rect 1593 5049 1627 5083
rect 2881 5049 2915 5083
rect 3801 5049 3835 5083
rect 1869 4981 1903 5015
rect 2145 4981 2179 5015
rect 2697 4981 2731 5015
rect 3617 4981 3651 5015
rect 5365 4981 5399 5015
rect 4629 4777 4663 4811
rect 4997 4777 5031 4811
rect 5365 4777 5399 4811
rect 5089 4641 5123 4675
rect 4445 4573 4479 4607
rect 4997 4573 5031 4607
rect 1593 4233 1627 4267
rect 1409 4097 1443 4131
rect 3525 4097 3559 4131
rect 3709 4097 3743 4131
rect 5181 4097 5215 4131
rect 3893 4029 3927 4063
rect 5365 3893 5399 3927
rect 2237 3689 2271 3723
rect 2053 3485 2087 3519
rect 2237 3485 2271 3519
rect 2789 3009 2823 3043
rect 2973 2805 3007 2839
rect 1869 2601 1903 2635
rect 3801 2601 3835 2635
rect 1593 2533 1627 2567
rect 4077 2465 4111 2499
rect 4169 2465 4203 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3985 2397 4019 2431
rect 4261 2397 4295 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 1394 8984 1400 9036
rect 1452 8984 1458 9036
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 3142 8956 3148 8968
rect 1719 8928 3148 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 842 8440 848 8492
rect 900 8480 906 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 900 8452 1409 8480
rect 900 8440 906 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 3050 8440 3056 8492
rect 3108 8480 3114 8492
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 3108 8452 3157 8480
rect 3108 8440 3114 8452
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3510 8480 3516 8492
rect 3375 8452 3516 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 3234 8344 3240 8356
rect 1627 8316 3240 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 4890 8344 4896 8356
rect 3375 8316 4896 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2958 7868 2964 7880
rect 2547 7840 2964 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2424 7800 2452 7831
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4672 7840 5181 7868
rect 4672 7828 4678 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5258 7800 5264 7812
rect 2424 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1762 7732 1768 7744
rect 1627 7704 1768 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 4338 7732 4344 7744
rect 2731 7704 4344 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 3234 7488 3240 7540
rect 3292 7488 3298 7540
rect 3252 7460 3280 7488
rect 3068 7432 3280 7460
rect 3068 7401 3096 7432
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7361 3111 7395
rect 3053 7355 3111 7361
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3292 7364 4077 7392
rect 3292 7352 3298 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 3142 7284 3148 7336
rect 3200 7284 3206 7336
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 3421 7259 3479 7265
rect 3421 7225 3433 7259
rect 3467 7256 3479 7259
rect 5166 7256 5172 7268
rect 3467 7228 5172 7256
rect 3467 7225 3479 7228
rect 3421 7219 3479 7225
rect 5166 7216 5172 7228
rect 5224 7216 5230 7268
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4982 7188 4988 7200
rect 4479 7160 4988 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4212 6752 4813 6780
rect 4212 6740 4218 6752
rect 4801 6749 4813 6752
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 1854 6712 1860 6724
rect 1596 6684 1860 6712
rect 1596 6653 1624 6684
rect 1854 6672 1860 6684
rect 1912 6712 1918 6724
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 1912 6684 5181 6712
rect 1912 6672 1918 6684
rect 5169 6681 5181 6684
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 5074 6604 5080 6656
rect 5132 6604 5138 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 2958 6400 2964 6452
rect 3016 6400 3022 6452
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3326 6304 3332 6316
rect 3283 6276 3332 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 5132 6276 5181 6304
rect 5132 6264 5138 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 1820 6208 2973 6236
rect 1820 6196 1826 6208
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3418 6100 3424 6112
rect 3200 6072 3424 6100
rect 3200 6060 3206 6072
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 3418 5352 3424 5364
rect 1688 5324 3424 5352
rect 1688 5293 1716 5324
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 4430 5352 4436 5364
rect 3559 5324 4436 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4798 5352 4804 5364
rect 4571 5324 4804 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5253 1731 5287
rect 3326 5284 3332 5296
rect 1673 5247 1731 5253
rect 1780 5256 3332 5284
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1780 5157 1808 5256
rect 3326 5244 3332 5256
rect 3384 5244 3390 5296
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1912 5188 1961 5216
rect 1912 5176 1918 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2648 5188 2697 5216
rect 2648 5176 2654 5188
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 3142 5176 3148 5228
rect 3200 5176 3206 5228
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 4341 5219 4399 5225
rect 4341 5216 4353 5219
rect 3476 5188 4353 5216
rect 3476 5176 3482 5188
rect 4341 5185 4353 5188
rect 4387 5216 4399 5219
rect 4522 5216 4528 5228
rect 4387 5188 4528 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4890 5176 4896 5228
rect 4948 5216 4954 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4948 5188 5181 5216
rect 4948 5176 4954 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2314 5108 2320 5160
rect 2372 5148 2378 5160
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2372 5120 2513 5148
rect 2372 5108 2378 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 3050 5108 3056 5160
rect 3108 5108 3114 5160
rect 4062 5108 4068 5160
rect 4120 5108 4126 5160
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5080 1639 5083
rect 2590 5080 2596 5092
rect 1627 5052 2596 5080
rect 1627 5049 1639 5052
rect 1581 5043 1639 5049
rect 2590 5040 2596 5052
rect 2648 5040 2654 5092
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5080 2927 5083
rect 3789 5083 3847 5089
rect 3789 5080 3801 5083
rect 2915 5052 3801 5080
rect 2915 5049 2927 5052
rect 2869 5043 2927 5049
rect 3789 5049 3801 5052
rect 3835 5080 3847 5083
rect 3970 5080 3976 5092
rect 3835 5052 3976 5080
rect 3835 5049 3847 5052
rect 3789 5043 3847 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 1854 4972 1860 5024
rect 1912 4972 1918 5024
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 2406 5012 2412 5024
rect 2179 4984 2412 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 2685 5015 2743 5021
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 3142 5012 3148 5024
rect 2731 4984 3148 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 3602 4972 3608 5024
rect 3660 4972 3666 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 4614 4768 4620 4820
rect 4672 4768 4678 4820
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4777 5043 4811
rect 4985 4771 5043 4777
rect 3326 4700 3332 4752
rect 3384 4740 3390 4752
rect 5000 4740 5028 4771
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 5316 4780 5365 4808
rect 5316 4768 5322 4780
rect 5353 4777 5365 4780
rect 5399 4777 5411 4811
rect 5353 4771 5411 4777
rect 3384 4712 5028 4740
rect 3384 4700 3390 4712
rect 1854 4632 1860 4684
rect 1912 4672 1918 4684
rect 5077 4675 5135 4681
rect 5077 4672 5089 4675
rect 1912 4644 5089 4672
rect 1912 4632 1918 4644
rect 5077 4641 5089 4644
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4396 4576 4445 4604
rect 4396 4564 4402 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4580 4576 4997 4604
rect 4580 4564 4586 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 1581 4267 1639 4273
rect 1581 4233 1593 4267
rect 1627 4264 1639 4267
rect 3142 4264 3148 4276
rect 1627 4236 3148 4264
rect 1627 4233 1639 4236
rect 1581 4227 1639 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4154 4128 4160 4140
rect 3743 4100 4160 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 3712 4060 3740 4091
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4488 4100 5181 4128
rect 4488 4088 4494 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 2464 4032 3740 4060
rect 3881 4063 3939 4069
rect 2464 4020 2470 4032
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 3970 4060 3976 4072
rect 3927 4032 3976 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 3050 3720 3056 3732
rect 2271 3692 3056 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 2498 3584 2504 3596
rect 2056 3556 2504 3584
rect 2056 3525 2084 3556
rect 2498 3544 2504 3556
rect 2556 3584 2562 3596
rect 3970 3584 3976 3596
rect 2556 3556 3976 3584
rect 2556 3544 2562 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2406 3516 2412 3528
rect 2271 3488 2412 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 3602 3040 3608 3052
rect 2823 3012 3608 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 4614 2836 4620 2848
rect 3007 2808 4620 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 3234 2632 3240 2644
rect 1903 2604 3240 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 4062 2632 4068 2644
rect 3835 2604 4068 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 2314 2564 2320 2576
rect 1627 2536 2320 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 2314 2524 2320 2536
rect 2372 2564 2378 2576
rect 2372 2536 4292 2564
rect 2372 2524 2378 2536
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3200 2468 4077 2496
rect 3200 2456 3206 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4154 2456 4160 2508
rect 4212 2456 4218 2508
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 4264 2437 4292 2536
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 5040 2400 5089 2428
rect 5040 2388 5046 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 3148 8916 3200 8968
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 848 8440 900 8492
rect 3056 8440 3108 8492
rect 3516 8440 3568 8492
rect 3240 8304 3292 8356
rect 4896 8304 4948 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 848 7828 900 7880
rect 2964 7828 3016 7880
rect 4620 7828 4672 7880
rect 5264 7760 5316 7812
rect 1768 7692 1820 7744
rect 4344 7692 4396 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 3240 7488 3292 7540
rect 3240 7352 3292 7404
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 5172 7216 5224 7268
rect 4988 7148 5040 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 848 6740 900 6792
rect 4160 6740 4212 6792
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 1860 6672 1912 6724
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 3332 6264 3384 6316
rect 5080 6264 5132 6316
rect 1768 6196 1820 6248
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 3424 6060 3476 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 3424 5312 3476 5364
rect 4436 5312 4488 5364
rect 4804 5312 4856 5364
rect 848 5176 900 5228
rect 3332 5244 3384 5296
rect 1860 5176 1912 5228
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2596 5176 2648 5228
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 3424 5176 3476 5228
rect 4528 5176 4580 5228
rect 4896 5176 4948 5228
rect 2320 5108 2372 5160
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 2596 5040 2648 5092
rect 3976 5040 4028 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2412 4972 2464 5024
rect 3148 4972 3200 5024
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 3332 4700 3384 4752
rect 5264 4768 5316 4820
rect 1860 4632 1912 4684
rect 4344 4564 4396 4616
rect 4528 4564 4580 4616
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 3148 4224 3200 4276
rect 848 4088 900 4140
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 2412 4020 2464 4072
rect 4160 4088 4212 4140
rect 4436 4088 4488 4140
rect 3976 4020 4028 4072
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 3056 3680 3108 3732
rect 2504 3544 2556 3596
rect 3976 3544 4028 3596
rect 2412 3476 2464 3528
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 3608 3000 3660 3052
rect 4620 2796 4672 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 3240 2592 3292 2644
rect 4068 2592 4120 2644
rect 2320 2524 2372 2576
rect 3148 2456 3200 2508
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 4160 2456 4212 2465
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 4988 2388 5040 2440
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 1412 9042 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 1400 9036 1452 9042
rect 5354 9007 5410 9016
rect 1400 8978 1452 8984
rect 3148 8968 3200 8974
rect 846 8936 902 8945
rect 3148 8910 3200 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 846 8871 902 8880
rect 860 8498 888 8871
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 848 7880 900 7886
rect 846 7848 848 7857
rect 2964 7880 3016 7886
rect 900 7848 902 7857
rect 2964 7822 3016 7828
rect 846 7783 902 7792
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 1780 6254 1808 7686
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 846 5128 902 5137
rect 1780 5114 1808 6190
rect 1872 5234 1900 6666
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2976 6458 3004 7822
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2320 5160 2372 5166
rect 1780 5086 1900 5114
rect 2320 5102 2372 5108
rect 846 5063 902 5072
rect 1872 5030 1900 5086
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 4690 1900 4966
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 3777 888 4082
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 846 3768 902 3777
rect 1950 3771 2258 3780
rect 846 3703 902 3712
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2332 2582 2360 5102
rect 2424 5030 2452 5170
rect 2608 5114 2636 5170
rect 3068 5166 3096 8434
rect 3160 7342 3188 8910
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 7562 3280 8298
rect 3252 7546 3372 7562
rect 3240 7540 3372 7546
rect 3292 7534 3372 7540
rect 3240 7482 3292 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3160 6118 3188 7278
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 2516 5098 2636 5114
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2516 5092 2648 5098
rect 2516 5086 2596 5092
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2424 4078 2452 4966
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2424 3534 2452 4014
rect 2516 3602 2544 5086
rect 2596 5034 2648 5040
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 3068 3738 3096 5102
rect 3160 5030 3188 5170
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3160 4282 3188 4966
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 3160 2514 3188 4218
rect 3252 2650 3280 7346
rect 3344 6322 3372 7534
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3344 5302 3372 6258
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5370 3464 6054
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3344 4758 3372 5238
rect 3436 5234 3464 5306
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3528 4146 3556 8434
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 5098 4016 7278
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3620 3058 3648 4966
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3988 3602 4016 4014
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3988 2446 4016 3538
rect 4080 2650 4108 5102
rect 4172 4146 4200 6734
rect 4356 4622 4384 7686
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4448 4146 4476 5306
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4540 4622 4568 5170
rect 4632 4826 4660 7822
rect 4816 5370 4844 8910
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4908 5234 4936 8298
rect 5184 7274 5212 8910
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4172 2514 4200 4082
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4632 2446 4660 2790
rect 5000 2446 5028 7142
rect 5276 6798 5304 7754
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6322 5120 6598
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5276 4826 5304 6734
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 6361 5396 6394
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 846 8880 902 8936
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 846 7828 848 7848
rect 848 7828 900 7848
rect 900 7828 902 7848
rect 846 7792 902 7828
rect 846 6432 902 6488
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 846 5072 902 5128
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 846 3712 902 3768
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5354 3576 5410 3632
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7850 907 7853
rect 798 7848 907 7850
rect 798 7792 846 7848
rect 902 7792 907 7848
rect 798 7787 907 7792
rect 798 7744 858 7787
rect 0 7654 858 7744
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 0 7624 800 7654
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__or4_2  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_
timestamp 1704896540
transform -1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _16_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp 1704896540
transform 1 0 2852 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 1704896540
transform 1 0 2300 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1704896540
transform -1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1704896540
transform -1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_21
timestamp 1704896540
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_33
timestamp 1704896540
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_45
timestamp 1704896540
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_9
timestamp 1704896540
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_13
timestamp 1704896540
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1704896540
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 1704896540
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 1704896540
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_31
timestamp 1704896540
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_43
timestamp 1704896540
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_35
timestamp 1704896540
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_39
timestamp 1704896540
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 1704896540
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_13
timestamp 1704896540
transform 1 0 2300 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_33
timestamp 1704896540
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_38
timestamp 1704896540
transform 1 0 4600 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 1704896540
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_19
timestamp 1704896540
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_24
timestamp 1704896540
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_36
timestamp 1704896540
transform 1 0 4416 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 1704896540
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1704896540
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_37
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_46
timestamp 1704896540
transform 1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_26
timestamp 1704896540
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_37
timestamp 1704896540
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_45
timestamp 1704896540
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_6
timestamp 1704896540
transform 1 0 1656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_12
timestamp 1704896540
transform 1 0 2208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1704896540
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1704896540
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_18
timestamp 1704896540
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_25
timestamp 1704896540
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_37
timestamp 1704896540
transform 1 0 4508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_45
timestamp 1704896540
transform 1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1704896540
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1704896540
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1704896540
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704896540
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 in[0]
port 2 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 in[1]
port 3 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 in[2]
port 4 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 in[3]
port 5 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 in[4]
port 6 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 in[5]
port 7 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 in[6]
port 8 nsew signal input
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 in[7]
port 9 nsew signal input
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 480 0 0 0 out[0]
port 10 nsew signal output
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 480 0 0 0 out[1]
port 11 nsew signal output
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 480 0 0 0 out[2]
port 12 nsew signal output
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 480 0 0 0 out[3]
port 13 nsew signal output
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 480 0 0 0 out[4]
port 14 nsew signal output
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 480 0 0 0 out[5]
port 15 nsew signal output
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 480 0 0 0 out[6]
port 16 nsew signal output
flabel metal3 s 6100 824 6900 944 0 FreeSans 480 0 0 0 out[7]
port 17 nsew signal output
rlabel metal1 3450 8704 3450 8704 0 VGND
rlabel metal1 3450 9248 3450 9248 0 VPWR
rlabel metal1 3956 4114 3956 4114 0 _00_
rlabel metal2 3082 4420 3082 4420 0 _01_
rlabel metal1 3450 8466 3450 8466 0 _02_
rlabel metal1 3956 2618 3956 2618 0 _03_
rlabel metal1 3910 5066 3910 5066 0 _04_
rlabel metal1 3220 3026 3220 3026 0 _05_
rlabel metal2 5290 5780 5290 5780 0 _06_
rlabel metal1 2760 7854 2760 7854 0 _07_
rlabel metal1 4416 4590 4416 4590 0 _08_
rlabel metal3 1050 10404 1050 10404 0 in[0]
rlabel metal3 751 9044 751 9044 0 in[1]
rlabel metal3 751 7684 751 7684 0 in[2]
rlabel metal3 751 6324 751 6324 0 in[3]
rlabel metal3 751 4964 751 4964 0 in[4]
rlabel metal3 751 3604 751 3604 0 in[5]
rlabel metal3 751 2244 751 2244 0 in[6]
rlabel metal3 1188 884 1188 884 0 in[7]
rlabel metal1 4462 5202 4462 5202 0 net1
rlabel metal1 4324 7242 4324 7242 0 net10
rlabel metal1 4922 7854 4922 7854 0 net11
rlabel metal1 5152 6290 5152 6290 0 net12
rlabel metal1 5060 5202 5060 5202 0 net13
rlabel metal1 4830 4114 4830 4114 0 net14
rlabel metal2 4646 2618 4646 2618 0 net15
rlabel metal1 5060 2414 5060 2414 0 net16
rlabel metal1 3312 6290 3312 6290 0 net2
rlabel metal2 1886 4828 1886 4828 0 net3
rlabel metal1 1610 6664 1610 6664 0 net4
rlabel metal1 3956 4046 3956 4046 0 net5
rlabel metal2 3174 3842 3174 3842 0 net6
rlabel metal1 2944 2550 2944 2550 0 net7
rlabel metal1 2576 2618 2576 2618 0 net8
rlabel metal1 4692 5338 4692 5338 0 net9
rlabel metal2 5014 9775 5014 9775 0 out[0]
rlabel via2 5382 9061 5382 9061 0 out[1]
rlabel via2 5382 7701 5382 7701 0 out[2]
rlabel metal2 5382 6375 5382 6375 0 out[3]
rlabel via2 5382 4981 5382 4981 0 out[4]
rlabel metal2 5382 3757 5382 3757 0 out[5]
rlabel via2 4830 2261 4830 2261 0 out[6]
rlabel metal2 5474 1615 5474 1615 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
