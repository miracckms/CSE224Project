magic
tech sky130A
magscale 1 2
timestamp 1745676756
<< checkpaint >>
rect -3932 -3108 10832 14396
<< viali >>
rect 2973 9129 3007 9163
rect 4997 9129 5031 9163
rect 5365 9061 5399 9095
rect 1409 8993 1443 9027
rect 1685 8925 1719 8959
rect 2881 8925 2915 8959
rect 2973 8925 3007 8959
rect 3801 8925 3835 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 3157 8857 3191 8891
rect 2697 8789 2731 8823
rect 4077 8789 4111 8823
rect 1593 8585 1627 8619
rect 1409 8449 1443 8483
rect 1593 8041 1627 8075
rect 4077 8041 4111 8075
rect 2237 7973 2271 8007
rect 3617 7905 3651 7939
rect 4261 7905 4295 7939
rect 1409 7837 1443 7871
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2421 7837 2455 7871
rect 2697 7837 2731 7871
rect 2881 7837 2915 7871
rect 3433 7837 3467 7871
rect 3985 7837 4019 7871
rect 5181 7837 5215 7871
rect 2605 7769 2639 7803
rect 2789 7701 2823 7735
rect 3249 7701 3283 7735
rect 4261 7701 4295 7735
rect 5365 7701 5399 7735
rect 4261 7497 4295 7531
rect 2329 7361 2363 7395
rect 3893 7361 3927 7395
rect 3985 7361 4019 7395
rect 2513 7225 2547 7259
rect 3893 7157 3927 7191
rect 1593 6885 1627 6919
rect 1409 6749 1443 6783
rect 2421 6749 2455 6783
rect 5181 6749 5215 6783
rect 2605 6613 2639 6647
rect 5365 6613 5399 6647
rect 3893 6273 3927 6307
rect 3985 6205 4019 6239
rect 4261 6205 4295 6239
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 2237 5525 2271 5559
rect 4813 5321 4847 5355
rect 1409 5185 1443 5219
rect 4997 5185 5031 5219
rect 5181 5185 5215 5219
rect 1593 4981 1627 5015
rect 5365 4981 5399 5015
rect 1409 4097 1443 4131
rect 3617 4097 3651 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 3525 4029 3559 4063
rect 1593 3961 1627 3995
rect 3985 3961 4019 3995
rect 4169 3961 4203 3995
rect 4077 3893 4111 3927
rect 5365 3893 5399 3927
rect 4629 3689 4663 3723
rect 4813 3485 4847 3519
rect 4905 3485 4939 3519
rect 4537 3145 4571 3179
rect 2789 3009 2823 3043
rect 4077 3009 4111 3043
rect 4261 3009 4295 3043
rect 4353 3009 4387 3043
rect 2881 2941 2915 2975
rect 3157 2805 3191 2839
rect 4077 2805 4111 2839
rect 1593 2601 1627 2635
rect 1869 2601 1903 2635
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 2958 9120 2964 9172
rect 3016 9120 3022 9172
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 1394 8984 1400 9036
rect 1452 8984 1458 9036
rect 3142 9024 3148 9036
rect 2884 8996 3148 9024
rect 2884 8965 2912 8996
rect 3142 8984 3148 8996
rect 3200 9024 3206 9036
rect 3200 8996 4200 9024
rect 3200 8984 3206 8996
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3050 8956 3056 8968
rect 3007 8928 3056 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 1688 8888 1716 8919
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 4172 8965 4200 8996
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4338 8956 4344 8968
rect 4295 8928 4344 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 3145 8891 3203 8897
rect 3145 8888 3157 8891
rect 1688 8860 3157 8888
rect 3145 8857 3157 8860
rect 3191 8888 3203 8891
rect 3694 8888 3700 8900
rect 3191 8860 3700 8888
rect 3191 8857 3203 8860
rect 3145 8851 3203 8857
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2556 8792 2697 8820
rect 2556 8780 2562 8792
rect 2685 8789 2697 8792
rect 2731 8820 2743 8823
rect 3804 8820 3832 8919
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 2731 8792 3832 8820
rect 2731 8789 2743 8792
rect 2685 8783 2743 8789
rect 4062 8780 4068 8832
rect 4120 8780 4126 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 3050 8616 3056 8628
rect 1627 8588 3056 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 3050 8576 3056 8588
rect 3108 8616 3114 8628
rect 3878 8616 3884 8628
rect 3108 8588 3884 8616
rect 3108 8576 3114 8588
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 842 8440 848 8492
rect 900 8480 906 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 900 8452 1409 8480
rect 900 8440 906 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2958 8072 2964 8084
rect 1627 8044 2964 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3694 8032 3700 8084
rect 3752 8072 3758 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3752 8044 4077 8072
rect 3752 8032 3758 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 2225 8007 2283 8013
rect 2225 7973 2237 8007
rect 2271 8004 2283 8007
rect 2498 8004 2504 8016
rect 2271 7976 2504 8004
rect 2271 7973 2283 7976
rect 2225 7967 2283 7973
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 2976 8004 3004 8032
rect 3970 8004 3976 8016
rect 2976 7976 3976 8004
rect 3970 7964 3976 7976
rect 4028 8004 4034 8016
rect 4028 7976 4292 8004
rect 4028 7964 4034 7976
rect 1578 7896 1584 7948
rect 1636 7936 1642 7948
rect 4264 7945 4292 7976
rect 3605 7939 3663 7945
rect 3605 7936 3617 7939
rect 1636 7908 2452 7936
rect 1636 7896 1642 7908
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 1728 7840 2145 7868
rect 1728 7828 1734 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 2424 7877 2452 7908
rect 2700 7908 3617 7936
rect 2700 7877 2728 7908
rect 3605 7905 3617 7908
rect 3651 7905 3663 7939
rect 3605 7899 3663 7905
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2455 7840 2697 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2832 7840 2881 7868
rect 2832 7828 2838 7840
rect 2869 7837 2881 7840
rect 2915 7868 2927 7871
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 2915 7840 3433 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3421 7837 3433 7840
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3878 7868 3884 7880
rect 3568 7840 3884 7868
rect 3568 7828 3574 7840
rect 3878 7828 3884 7840
rect 3936 7868 3942 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3936 7840 3985 7868
rect 3936 7828 3942 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4212 7840 5181 7868
rect 4212 7828 4218 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 2593 7803 2651 7809
rect 2593 7769 2605 7803
rect 2639 7800 2651 7803
rect 4522 7800 4528 7812
rect 2639 7772 4528 7800
rect 2639 7769 2651 7772
rect 2593 7763 2651 7769
rect 4522 7760 4528 7772
rect 4580 7760 4586 7812
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 2958 7732 2964 7744
rect 2823 7704 2964 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3234 7692 3240 7744
rect 3292 7692 3298 7744
rect 4246 7692 4252 7744
rect 4304 7692 4310 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4338 7528 4344 7540
rect 4295 7500 4344 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4338 7488 4344 7500
rect 4396 7528 4402 7540
rect 4890 7528 4896 7540
rect 4396 7500 4896 7528
rect 4396 7488 4402 7500
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 3694 7420 3700 7472
rect 3752 7460 3758 7472
rect 3752 7432 3924 7460
rect 3752 7420 3758 7432
rect 3896 7404 3924 7432
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 3786 7392 3792 7404
rect 2363 7364 3792 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 3878 7352 3884 7404
rect 3936 7352 3942 7404
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7256 2559 7259
rect 4430 7256 4436 7268
rect 2547 7228 4436 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 4430 7216 4436 7228
rect 4488 7216 4494 7268
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3568 7160 3893 7188
rect 3568 7148 3574 7160
rect 3881 7157 3893 7160
rect 3927 7188 3939 7191
rect 3970 7188 3976 7200
rect 3927 7160 3976 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 1581 6919 1639 6925
rect 1581 6885 1593 6919
rect 1627 6914 1639 6919
rect 1627 6886 1661 6914
rect 1627 6885 1639 6886
rect 1581 6879 1639 6885
rect 1596 6848 1624 6879
rect 3142 6848 3148 6860
rect 1596 6820 3148 6848
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 2424 6712 2452 6743
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 4120 6752 5181 6780
rect 4120 6740 4126 6752
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 4614 6712 4620 6724
rect 2424 6684 4620 6712
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 2593 6647 2651 6653
rect 2593 6613 2605 6647
rect 2639 6644 2651 6647
rect 4154 6644 4160 6656
rect 2639 6616 4160 6644
rect 2639 6613 2651 6616
rect 2593 6607 2651 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 3988 6304 4016 6332
rect 3927 6276 4016 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 3970 6196 3976 6248
rect 4028 6196 4034 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 5166 6236 5172 6248
rect 4295 6208 5172 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 3234 5692 3240 5704
rect 2363 5664 3240 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2148 5624 2176 5655
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 2958 5624 2964 5636
rect 2148 5596 2964 5624
rect 2958 5584 2964 5596
rect 3016 5624 3022 5636
rect 3510 5624 3516 5636
rect 3016 5596 3516 5624
rect 3016 5584 3022 5596
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 5166 5556 5172 5568
rect 2271 5528 5172 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 4798 5312 4804 5364
rect 4856 5312 4862 5364
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4028 5188 4997 5216
rect 4028 5176 4034 5188
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5166 5176 5172 5228
rect 5224 5176 5230 5228
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 2372 4100 3617 4128
rect 2372 4088 2378 4100
rect 3605 4097 3617 4100
rect 3651 4128 3663 4131
rect 4062 4128 4068 4140
rect 3651 4100 4068 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 3510 4020 3516 4072
rect 3568 4020 3574 4072
rect 5184 4060 5212 4091
rect 3988 4032 5212 4060
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2314 3992 2320 4004
rect 1627 3964 2320 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2314 3952 2320 3964
rect 2372 3952 2378 4004
rect 3988 4001 4016 4032
rect 3973 3995 4031 4001
rect 3973 3961 3985 3995
rect 4019 3961 4031 3995
rect 3973 3955 4031 3961
rect 4154 3952 4160 4004
rect 4212 3952 4218 4004
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3844 3896 4077 3924
rect 3844 3884 3850 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 4614 3680 4620 3732
rect 4672 3680 4678 3732
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4304 3488 4813 3516
rect 4304 3476 4310 3488
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 1578 3340 1584 3392
rect 1636 3380 1642 3392
rect 4338 3380 4344 3392
rect 1636 3352 4344 3380
rect 1636 3340 1642 3352
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 4154 3176 4160 3188
rect 2924 3148 4160 3176
rect 2924 3136 2930 3148
rect 4154 3136 4160 3148
rect 4212 3176 4218 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4212 3148 4537 3176
rect 4212 3136 4218 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 1728 3080 4292 3108
rect 1728 3068 1734 3080
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 4264 3049 4292 3080
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 3160 3012 4077 3040
rect 2866 2932 2872 2984
rect 2924 2932 2930 2984
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 3160 2904 3188 3012
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 5074 2904 5080 2916
rect 2556 2876 3188 2904
rect 3252 2876 5080 2904
rect 2556 2864 2562 2876
rect 3145 2839 3203 2845
rect 3145 2805 3157 2839
rect 3191 2836 3203 2839
rect 3252 2836 3280 2876
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 3191 2808 3280 2836
rect 3191 2805 3203 2808
rect 3145 2799 3203 2805
rect 4062 2796 4068 2848
rect 4120 2796 4126 2848
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 1670 2632 1676 2644
rect 1627 2604 1676 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2774 2632 2780 2644
rect 1903 2604 2780 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4488 2400 4629 2428
rect 4488 2388 4494 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 3148 8984 3200 9036
rect 3056 8916 3108 8968
rect 3700 8848 3752 8900
rect 2504 8780 2556 8832
rect 4344 8916 4396 8968
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 4068 8823 4120 8832
rect 4068 8789 4077 8823
rect 4077 8789 4111 8823
rect 4111 8789 4120 8823
rect 4068 8780 4120 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 3056 8576 3108 8628
rect 3884 8576 3936 8628
rect 848 8440 900 8492
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 2964 8032 3016 8084
rect 3700 8032 3752 8084
rect 2504 7964 2556 8016
rect 3976 7964 4028 8016
rect 1584 7896 1636 7948
rect 848 7828 900 7880
rect 1676 7828 1728 7880
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 2780 7828 2832 7880
rect 3516 7828 3568 7880
rect 3884 7828 3936 7880
rect 4160 7828 4212 7880
rect 4528 7760 4580 7812
rect 2964 7692 3016 7744
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 4344 7488 4396 7540
rect 4896 7488 4948 7540
rect 3700 7420 3752 7472
rect 3792 7352 3844 7404
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4436 7216 4488 7268
rect 3516 7148 3568 7200
rect 3976 7148 4028 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 3148 6808 3200 6860
rect 848 6740 900 6792
rect 4068 6740 4120 6792
rect 4620 6672 4672 6724
rect 4160 6604 4212 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 3976 6332 4028 6384
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 5172 6196 5224 6248
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 3240 5652 3292 5704
rect 2964 5584 3016 5636
rect 3516 5584 3568 5636
rect 5172 5516 5224 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 4804 5355 4856 5364
rect 4804 5321 4813 5355
rect 4813 5321 4847 5355
rect 4847 5321 4856 5355
rect 4804 5312 4856 5321
rect 848 5176 900 5228
rect 3976 5176 4028 5228
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 848 4088 900 4140
rect 2320 4088 2372 4140
rect 4068 4088 4120 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 3516 4063 3568 4072
rect 3516 4029 3525 4063
rect 3525 4029 3559 4063
rect 3559 4029 3568 4063
rect 3516 4020 3568 4029
rect 2320 3952 2372 4004
rect 4160 3995 4212 4004
rect 4160 3961 4169 3995
rect 4169 3961 4203 3995
rect 4203 3961 4212 3995
rect 4160 3952 4212 3961
rect 3792 3884 3844 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 4252 3476 4304 3528
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 1584 3340 1636 3392
rect 4344 3340 4396 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 2872 3136 2924 3188
rect 4160 3136 4212 3188
rect 1676 3068 1728 3120
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 2504 2864 2556 2916
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 5080 2864 5132 2916
rect 4068 2839 4120 2848
rect 4068 2805 4077 2839
rect 4077 2805 4111 2839
rect 4111 2805 4120 2839
rect 4068 2796 4120 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 1676 2592 1728 2644
rect 2780 2592 2832 2644
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4436 2388 4488 2440
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 1412 9042 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 846 8936 902 8945
rect 846 8871 902 8880
rect 860 8498 888 8871
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2516 8022 2544 8774
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2976 8090 3004 9114
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 3148 9036 3200 9042
rect 5354 9007 5410 9016
rect 3148 8978 3200 8984
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8634 3096 8910
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 848 7880 900 7886
rect 846 7848 848 7857
rect 900 7848 902 7857
rect 846 7783 902 7792
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 846 5128 902 5137
rect 846 5063 902 5072
rect 1596 5030 1624 7890
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2516 7834 2544 7958
rect 2780 7880 2832 7886
rect 2516 7828 2780 7834
rect 2516 7822 2832 7828
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 3777 888 4082
rect 846 3768 902 3777
rect 846 3703 902 3712
rect 1596 3398 1624 4966
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1688 3126 1716 7822
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2332 4146 2360 7822
rect 2516 7806 2820 7822
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2332 4010 2360 4082
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1688 2650 1716 3062
rect 2516 2922 2544 7806
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2976 5642 3004 7686
rect 3160 6866 3188 8978
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3712 8090 3740 8842
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3252 5710 3280 7686
rect 3528 7206 3556 7822
rect 3712 7478 3740 8026
rect 3896 7886 3924 8570
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 3988 7410 4016 7958
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 3528 4078 3556 5578
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3804 3942 3832 7346
rect 3896 6202 3924 7346
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6390 4016 7142
rect 4080 6798 4108 8774
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4172 6662 4200 7822
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3976 6248 4028 6254
rect 3896 6196 3976 6202
rect 3896 6190 4028 6196
rect 3896 6174 4016 6190
rect 3988 5234 4016 6174
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2792 2650 2820 2994
rect 2884 2990 2912 3130
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 4080 2854 4108 4082
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3194 4200 3946
rect 4264 3534 4292 7686
rect 4356 7546 4384 8910
rect 4528 7812 4580 7818
rect 4528 7754 4580 7760
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4356 3058 4384 3334
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 4448 2446 4476 7210
rect 4540 4146 4568 7754
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4632 3738 4660 6666
rect 4816 5370 4844 8910
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4908 3534 4936 7482
rect 5184 6254 5212 8910
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6361 5396 6598
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 5234 5212 5510
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5092 2446 5120 2858
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 846 8880 902 8936
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 846 7828 848 7848
rect 848 7828 900 7848
rect 900 7828 902 7848
rect 846 7792 902 7828
rect 846 6432 902 6488
rect 846 5072 902 5128
rect 846 3712 902 3768
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5354 3576 5410 3632
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7850 907 7853
rect 798 7848 907 7850
rect 798 7792 846 7848
rect 902 7792 907 7848
rect 798 7787 907 7792
rect 798 7744 858 7787
rect 0 7654 858 7744
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 0 7624 800 7654
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__or4_2  _09_
timestamp 0
transform -1 0 3220 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_
timestamp 0
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_
timestamp 0
transform -1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _13_
timestamp 0
transform 1 0 3404 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _14_
timestamp 0
transform -1 0 2668 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _15_
timestamp 0
transform 1 0 4048 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _16_
timestamp 0
transform -1 0 4600 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 0
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _18_
timestamp 0
transform 1 0 2576 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp 0
transform 1 0 3680 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _20_
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _21_
timestamp 0
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform -1 0 5060 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform -1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _24_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 0
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_23
timestamp 0
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_31
timestamp 0
transform 1 0 3956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_38
timestamp 0
transform 1 0 4600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_46
timestamp 0
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 0
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_43
timestamp 0
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 0
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_18
timestamp 0
transform 1 0 2760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_24
timestamp 0
transform 1 0 3312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_38
timestamp 0
transform 1 0 4600 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 0
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_30
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_38
timestamp 0
transform 1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_14
timestamp 0
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_35
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 0
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_6
timestamp 0
transform 1 0 1656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_17
timestamp 0
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_11
timestamp 0
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_16
timestamp 0
transform 1 0 2576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_28
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_35
timestamp 0
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 0
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_20
timestamp 0
transform 1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_35
timestamp 0
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_43
timestamp 0
transform 1 0 5060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 0
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 0
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_42
timestamp 0
transform 1 0 4968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_13
timestamp 0
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_35
timestamp 0
transform 1 0 4324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_39
timestamp 0
transform 1 0 4692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal1 s 2852 2890 2852 2890 4 _00_
rlabel metal1 s 2162 5644 2162 5644 4 _01_
rlabel metal1 s 2806 5678 2806 5678 4 _02_
rlabel metal1 s 3588 7786 3588 7786 4 _03_
rlabel metal1 s 3726 3162 3726 3162 4 _04_
rlabel metal1 s 3956 3910 3956 3910 4 _05_
rlabel metal1 s 4324 7514 4324 7514 4 _06_
rlabel metal1 s 4554 3502 4554 3502 4 _07_
rlabel metal2 s 4646 5202 4646 5202 4 _08_
rlabel metal3 s 1050 10404 1050 10404 4 in[0]
rlabel metal3 s 0 8984 800 9104 4 in[1]
port 4 nsew
rlabel metal3 s 0 7624 800 7744 4 in[2]
port 5 nsew
rlabel metal3 s 0 6264 800 6384 4 in[3]
port 6 nsew
rlabel metal3 s 0 4904 800 5024 4 in[4]
port 7 nsew
rlabel metal3 s 0 3544 800 3664 4 in[5]
port 8 nsew
rlabel metal3 s 0 2184 800 2304 4 in[6]
port 9 nsew
rlabel metal3 s 1188 884 1188 884 4 in[7]
rlabel metal2 s 4002 5712 4002 5712 4 net1
rlabel metal1 s 4738 6222 4738 6222 4 net10
rlabel metal1 s 3404 6630 3404 6630 4 net11
rlabel metal1 s 4646 6766 4646 6766 4 net12
rlabel metal2 s 5198 5372 5198 5372 4 net13
rlabel metal1 s 5198 4080 5198 4080 4 net14
rlabel metal1 s 4554 2414 4554 2414 4 net15
rlabel metal2 s 5106 2652 5106 2652 4 net16
rlabel metal1 s 4002 6324 4002 6324 4 net2
rlabel metal2 s 2990 8602 2990 8602 4 net3
rlabel metal1 s 2392 6834 2392 6834 4 net4
rlabel metal2 s 1610 4182 1610 4182 4 net5
rlabel metal1 s 1978 3978 1978 3978 4 net6
rlabel metal1 s 1656 2618 1656 2618 4 net7
rlabel metal1 s 2346 2618 2346 2618 4 net8
rlabel metal2 s 4830 7140 4830 7140 4 net9
rlabel metal2 s 5014 9775 5014 9775 4 out[0]
rlabel metal3 s 5382 9061 5382 9061 4 out[1]
rlabel metal3 s 5382 7701 5382 7701 4 out[2]
rlabel metal2 s 5382 6477 5382 6477 4 out[3]
rlabel metal3 s 5382 4981 5382 4981 4 out[4]
rlabel metal2 s 5382 3757 5382 3757 4 out[5]
rlabel metal3 s 4830 2261 4830 2261 4 out[6]
rlabel metal2 s 5474 1615 5474 1615 4 out[7]
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 10344 800 10464 0 FreeSans 600 0 0 0 in[0]
port 3 nsew
flabel metal3 s 400 9044 400 9044 0 FreeSans 600 0 0 0 in[1]
flabel metal3 s 400 7684 400 7684 0 FreeSans 600 0 0 0 in[2]
flabel metal3 s 400 6324 400 6324 0 FreeSans 600 0 0 0 in[3]
flabel metal3 s 400 4964 400 4964 0 FreeSans 600 0 0 0 in[4]
flabel metal3 s 400 3604 400 3604 0 FreeSans 600 0 0 0 in[5]
flabel metal3 s 400 2244 400 2244 0 FreeSans 600 0 0 0 in[6]
flabel metal3 s 0 824 800 944 0 FreeSans 600 0 0 0 in[7]
port 10 nsew
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 600 0 0 0 out[0]
port 11 nsew
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 600 0 0 0 out[2]
port 13 nsew
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 600 0 0 0 out[3]
port 14 nsew
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 600 0 0 0 out[4]
port 15 nsew
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 600 0 0 0 out[5]
port 16 nsew
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 6100 824 6900 944 0 FreeSans 600 0 0 0 out[7]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
